/*************************************************************************
   Copyright 2008 Ray Salemi

   Licensed under the Apache License, Version 2.0 (the "License");
   you may not use this file except in compliance with the License.
   You may obtain a copy of the License at

       http://www.apache.org/licenses/LICENSE-2.0

   Unless required by applicable law or agreed to in writing, software
   distributed under the License is distributed on an "AS IS" BASIS,
   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
   See the License for the specific language governing permissions and
   limitations under the License.
**************************************************************************/
//
// Module tiny_cache_lib.cpubus_sm.fsm
//
// Created:
//          by - rsalemi.UNKNOWN (MAW-RSALEMI-LT)
//          at - 15:17:22 11/ 1/2006
//
// Generated by Mentor Graphics' HDL Designer(TM) 2006.1 (Build 56) Beta
//
module cpubus_sm( 
   clk, 
   cpuwait, 
   go, 
   rst, 
   transaction_req, 
   cpu_rd, 
   cpu_wr, 
   done, 
   reset
);


// Internal Declarations

input        clk;
input        cpuwait;
input        go;
input        rst;
input  [1:0] transaction_req;
output       cpu_rd;
output       cpu_wr;
output       done;
output       reset;


wire clk;
wire cpuwait;
wire go;
wire rst;
wire [1:0] transaction_req;
reg cpu_rd;
reg cpu_wr;
reg done;
reg reset;
// Module Declarations
parameter NOTHING = 0;
parameter READ = 1;
parameter WRITE = 2;
parameter RESET = 3;

// State encoding
parameter 
          INIT    = 3'd0,
          DOREAD  = 3'd1,
          DOWRITE = 3'd2,
          DORESET = 3'd3,
          WRITE2  = 3'd4;

reg [2:0] current_state, next_state;
// pragma state_vector current_state

//-----------------------------------------------------------------
// Next State Block for machine csm
//-----------------------------------------------------------------
always @(
   cpuwait or 
   current_state or 
   go or 
   transaction_req
)
begin : next_state_block_proc
   case (current_state) 
      INIT: begin
         if (go == 0)
            next_state = INIT;
         else if (transaction_req == READ)
            next_state = DOREAD;
         else if (transaction_req == WRITE)
            next_state = DOWRITE;
         else if ( transaction_req == RESET)
            next_state = DORESET;
      end
      DOREAD: begin
         if (cpuwait == 1)
            next_state = DOREAD;
         else if (cpuwait == 0)
            next_state = INIT;
      end
      DOWRITE: begin
         next_state = WRITE2;
      end
      DORESET: begin
         next_state = INIT;
      end
      WRITE2: begin
         next_state = INIT;
      end
      default: 
         next_state = INIT;
   endcase
end // Next State Block

//-----------------------------------------------------------------
// Output Block for machine csm
//-----------------------------------------------------------------
always @(
   current_state
)
begin : output_block_proc
   // Default Assignment
   cpu_rd = 0;
   cpu_wr = 0;
   done = 1;
   reset = 0;

   // Combined Actions
   case (current_state) 
      DOREAD: begin
          cpu_rd = 1;
         done = 0;
      end
      DOWRITE: begin
         cpu_wr = 1;
         done = 0;
      end
      DORESET: begin
          reset = 1;
         done = 0;
      end
      WRITE2: begin
          cpu_wr = 1;
         done = 0;
      end
      default: begin
      end
   endcase
end // Output Block

//-----------------------------------------------------------------
// Clocked Block for machine csm
//-----------------------------------------------------------------
always @(
   posedge clk or 
   negedge rst
) 
begin : clocked_block_proc
   if (!rst) begin
      current_state <= INIT;
   end
   else 
   begin
      current_state <= next_state;
   end
end // Clocked Block

endmodule // cpubus_sm
