/*************************************************************************
   Copyright 2008 Ray Salemi

   Licensed under the Apache License, Version 2.0 (the "License");
   you may not use this file except in compliance with the License.
   You may obtain a copy of the License at

       http://www.apache.org/licenses/LICENSE-2.0

   Unless required by applicable law or agreed to in writing, software
   distributed under the License is distributed on an "AS IS" BASIS,
   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
   See the License for the specific language governing permissions and
   limitations under the License.
**************************************************************************/
//
// Module ch2.top.struct
//
// Created:
//          by - Ray.UNKNOWN (OFFICE)
//          at - 11:34:42 07/28/2007
//
// Generated by Mentor Graphics' HDL Designer(TM) 2006.1 (Build 72)
//


module top;

// Internal Declarations



// Local declarations

// Internal signal declarations
// Internal Declarations




// Local declarations

// Internal signal declarations
wire       active;
reg        clk;
wire       cpu_rd;
wire       cpu_wr;
wire [7:0] cpubus_address;
wire [7:0] cpubus_data;
wire       cpuwait;
wire [7:0] memory_address;
wire [7:0] memory_data;
wire       memory_rd;
wire       memory_wr;
wire       reset;
wire       response;
wire [2:0] trans;



// Instances
//  Instances
cpubus_monitor_sm cpubus_monitor(
   .clk            (clk),
   .cpu_data       (cpubus_data),
   .cpu_rd         (cpu_rd),
   .cpu_wr         (cpu_wr),
   .cpubus_address (cpubus_address),
   .cpuwait        (cpuwait),
   .reset          (reset),
   .active         (active),
   .response       (response),
   .trans          (trans)
);

memory main_mem(
   .clk            (clk),
   .memory_address (memory_address),
   .memory_rd      (memory_rd),
   .memory_wr      (memory_wr),
   .memory_data    (memory_data)
);

scoreboard #(0,1,2,3,4,5,6,7,1,2) design_checker(
   .active         (active),
   .clk            (clk),
   .cpu_rd         (cpu_rd),
   .cpu_wr         (cpu_wr),
   .cpubus_address (cpubus_address),
   .cpubus_data    (cpubus_data),
   .memory_address (memory_address),
   .memory_data    (memory_data),
   .memory_rd      (memory_rd),
   .memory_wr      (memory_wr),
   .reset          (reset),
   .response       (response),
   .trans          (trans)
);

tester test_runner(
   .clk            (clk),
   .cpuwait        (cpuwait),
   .cpu_rd         (cpu_rd),
   .cpu_wr         (cpu_wr),
   .cpubus_address (cpubus_address),
   .reset          (reset),
   .cpu_data       (cpubus_data)
);

tiny_cache_vhd DUT(
   .clk         (clk),
   .cpu_address (cpubus_address),
   .cpu_rd      (cpu_rd),
   .cpu_wr      (cpu_wr),
   .rst         (reset),
   .cpuwait     (cpuwait),
   .mem_address (memory_address),
   .mem_rd      (memory_rd),
   .mem_wr      (memory_wr),
   .cpu_data    (cpubus_data),
   .mem_data    (memory_data)
);

// HDL Embedded Text Block eb1
//
// HDL Embedded Text Block 1 eb1
// eb1 1                       

initial clk = 0;
//
// HDL Embedded Text Block eb2
//
always #10 clk = ~clk;
//

endmodule // top
// tiny_cache_tb
