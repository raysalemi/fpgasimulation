-- *******************************************************************
-- Copyright 2008 Ray Salemi

-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License. 
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- ********************************************************************
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.STD_LOGIC_UNSIGNED.all;

ENTITY threebitcounter IS
   PORT( 
      clk      : IN     std_logic;
      data_in  : IN     std_logic_vector ( 2 DOWNTO 0 );
      inc      : IN     std_logic;
      ld       : IN     std_logic;
      rst      : IN     std_logic;
      data_out : BUFFER std_logic_vector ( 2 DOWNTO 0 )
   );

-- Declarations

END threebitcounter ;

--
-- VHDL Architecture vhdl_assert.threebitcounter.flow
--
-- Created:
--          by - Ray.UNKNOWN (OFFICE)
--          at - 15:24:22 08/11/2007
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2006.1 (Build 72)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
ARCHITECTURE flow OF threebitcounter IS

BEGIN

   process0_proc : PROCESS (clk)
		BEGIN
			IF (clk'EVENT AND clk = '1') THEN
		 -- Synchronous Reset
		 IF (rst = '1') THEN
			  data_out <= "000" ;
		 ELSE
			 IF ld = '1' THEN
				 data_out <= data_in;
			 ELSIF inc = '1' THEN
				 -- synthesis translate_off
				 assert (data_out /= "111")
				 	report "Oi! Counter Overflow"
				 	severity warning;
				 -- synthesis translate_on
				 data_out <= std_logic_vector(data_out + "001");
			 END IF;
		 END IF;
			END IF;
	END PROCESS process0_proc;


END flow;
