/*************************************************************************
   Copyright 2008 Ray Salemi

   Licensed under the Apache License, Version 2.0 (the "License");
   you may not use this file except in compliance with the License.
   You may obtain a copy of the License at

       http://www.apache.org/licenses/LICENSE-2.0

   Unless required by applicable law or agreed to in writing, software
   distributed under the License is distributed on an "AS IS" BASIS,
   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
   See the License for the specific language governing permissions and
   limitations under the License.
**************************************************************************/
//
// Module tinyCache_lib.tiny_cache.struct
//
// Created:
//          by - rsalemi.UNKNOWN (MAW-RSALEMI-LT)
//          at - 08:08:35 05/11/2005
//
// Generated by Mentor Graphics' HDL Designer(TM) 2005.1 (Build 83)
//


module tiny_cache_vlog( 
   clk, 
   cpu_address, 
   cpu_rd, 
   cpu_wr, 
   reset, 
   cpuwait, 
   memory_address, 
   memory_rd, 
   memory_wr, 
   cpu_data, 
   memory_data
);


parameter CACHE_DEPTH = 16;
parameter DATA_WIDTH = 8;
parameter ADDRESS_WIDTH = 8;
// Non hierarchical state machine declarations
// State encoding
parameter HIT = 2'd0;
parameter WRITE = 2'd1;
parameter MISS = 2'd2;
parameter RESET = 2'd3;

// Internal Declarations

input        clk;
input  [7:0] cpu_address;
input        cpu_rd;
input        cpu_wr;
input        reset;
output       cpuwait;
output [7:0] memory_address;
output       memory_rd;
output       memory_wr;
inout  [7:0] cpu_data;
inout  [7:0] memory_data;


wire clk;
wire [7:0] cpu_address;
wire cpu_rd;
wire cpu_wr;
wire reset;
wire cpuwait;
wire [7:0] memory_address;
reg memory_rd;
reg memory_wr;
wire [7:0] cpu_data;
wire [7:0] memory_data;
reg [1:0] cache_control_current_state, cache_control_next_state;
// pragma state_vector cache_control_current_state


// Internal signal declarations
wire [3:0] cache_address;


reg [DATA_WIDTH-1 : 0] cache_ram [0 : CACHE_DEPTH - 1];
reg [ADDRESS_WIDTH-1:0]  key_ram [0 : CACHE_DEPTH - 1];
reg [CACHE_DEPTH-1 : 0] invalid ;

// Instances 
// HDL Embedded Text Block 1 data_buffers
// eb1 1    

assign cpu_data  = (cpu_rd) ? cache_ram[cache_address] : 8'HZZ;
assign memory_data = (memory_wr) ? cpu_data : 8'HZZ;
assign cache_address = cpu_address[3:0];
assign memory_address = cpu_address;   
assign cpuwait =  ((key_ram[cache_address] != cpu_address) ||
                           (invalid [cache_address]) )&& cpu_rd; 
// (cpu_wr && (cache_address == 1)) ||
                           
// HDL Embedded Block 2 cache_sm
// Non hierarchical state machine
//-----------------------------------------------------------------
// Next State Block for machine cache_control
//-----------------------------------------------------------------
always @(
   cache_control_current_state or 
   cpu_wr or 
   cpuwait
)
begin : cache_control_next_state_block_proc
   case (cache_control_current_state) 
      HIT: begin
         if (cpuwait)
            cache_control_next_state = MISS;
         else if (cpu_wr)
            cache_control_next_state = WRITE;
         else
            cache_control_next_state = HIT;
      end
      WRITE: begin
         cache_control_next_state = HIT;
      end
      MISS: begin
         cache_control_next_state = HIT;
      end
      RESET: begin
         cache_control_next_state = HIT;
      end
      default: 
         cache_control_next_state = RESET;
   endcase
end // Next State Block

//-----------------------------------------------------------------
// Output Block for machine cache_control
//-----------------------------------------------------------------
always @(
   cache_control_current_state
)
begin : cache_control_output_block_proc
   // Default Assignment
   memory_rd = 0;
   memory_wr = 0;

   // Combined Actions
   case (cache_control_current_state) 
      HIT: begin
         memory_wr = 0;
      end
      WRITE: begin
         memory_wr = 1;
      end
      MISS: begin
         memory_rd = 1;
      end
      default: begin
      end
   endcase
end // Output Block

//-----------------------------------------------------------------
// Clocked Block for machine cache_control
//-----------------------------------------------------------------
always @(
   posedge clk
) 
begin : cache_control_clocked_block_proc
   if (reset) begin
      cache_control_current_state = RESET;
   end
   else 
   begin
      case (cache_control_current_state) 
        
            WRITE: begin
               key_ram[cache_address] = cpu_address;
               invalid[cache_address] = 0;
               cache_ram[cache_address] = cpu_data;
            end
            MISS: begin
               cache_ram[cache_address] = memory_data;
               key_ram[cache_address] = cpu_address;
               invalid[cache_address] = 0;
            end
            RESET : begin
               invalid = 16'hFFFF;
            end
      endcase
      cache_control_current_state = cache_control_next_state;
   end
end // Clocked Block







endmodule // tiny_cache_vlog

