// Accellera Standard V2.3 Open Verification Library (OVL).
// Accellera Copyright (c) 2005-2008. All rights reserved.

`include "std_ovl_defines.h"

`module ovl_arbiter (clock, reset, enable, reqs, priorities, gnts, fire);

  parameter severity_level      = `OVL_SEVERITY_DEFAULT;
  parameter width               = 2;
  parameter priority_width      = 1;
  parameter min_cks             = 1;
  parameter max_cks             = 0;
  parameter one_cycle_gnt_check = 1;
  parameter priority_check      = 0;
  parameter arbitration_rule    = 0;
  parameter property_type       = `OVL_PROPERTY_DEFAULT;
  parameter msg                 = `OVL_MSG_DEFAULT;
  parameter coverage_level      = `OVL_COVER_DEFAULT;

  parameter clock_edge          = `OVL_CLOCK_EDGE_DEFAULT;
  parameter reset_polarity      = `OVL_RESET_POLARITY_DEFAULT;
  parameter gating_type         = `OVL_GATING_TYPE_DEFAULT;

  input                    clock, reset, enable;
  input  [width-1 : 0]     reqs;
  input  [width-1 : 0]     gnts;
  input  [(width*priority_width)-1 : 0] priorities;
  output [`OVL_FIRE_WIDTH-1 : 0]   fire;

  // Parameters that should not be edited
  parameter assert_name = "OVL_ARBITER";

  `include "std_ovl_reset.h"
  `include "std_ovl_clock.h"
  `include "std_ovl_cover.h"
  `include "std_ovl_task.h"
  `include "std_ovl_init.h"

`ifdef OVL_SVA
  `include "./sva05/ovl_arbiter_logic.sv"
  assign fire = {`OVL_FIRE_WIDTH{1'b0}}; // Tied low in V2.3
`endif

`endmodule // ovl_arbiter

